////////////////////////////////////////////////////////////////////////////////
// Copyright (c) 2009  Bluespec, Inc.   ALL RIGHTS RESERVED.
////////////////////////////////////////////////////////////////////////////////
//  Filename      : BusRange.bsv
//  Description   :
////////////////////////////////////////////////////////////////////////////////
package BusRange;

// Notes :

////////////////////////////////////////////////////////////////////////////////
/// Imports
////////////////////////////////////////////////////////////////////////////////
import DefaultValue      ::*;

////////////////////////////////////////////////////////////////////////////////
/// Types
////////////////////////////////////////////////////////////////////////////////
typedef struct {
   addr_t      base;
   addr_t      high;
   } AddressRange#(type addr_t) deriving (Bits, Eq);

instance DefaultValue#(AddressRange#(addr_t))
   provisos(Bits#(addr_t, s0));
   defaultValue = AddressRange {
      base: unpack('1),
      high: unpack(0)
      };
endinstance

typedef function Bool f(addr_t x) MatchAddr#(type addr_t);

////////////////////////////////////////////////////////////////////////////////
/// Functions
////////////////////////////////////////////////////////////////////////////////
function MatchAddr#(addr_t) addAddressRangeMatch(AddressRange#(addr_t) r)
   provisos( Bits#(addr_t, s0)
           , Ord#(addr_t)
           );
   function f(x);
      return ((x >= r.base) && (x <= r.high));
   endfunction
   return f;
endfunction

endpackage: BusRange

